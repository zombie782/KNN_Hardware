`ifndef _defs_sv_
`define _defs_sv_

	localparam REF_DATA_POINTS=100;
	localparam QUERY_DATA_POINTS=20;
	
	localparam QUERY_FILE="query.txt";
	localparam REF_FILE="ref.txt";
	
	localparam DATA_DIM=30;
	localparam DIM_PREC=12;
	localparam CLASSIFICATIONS=2;
	
	localparam K=19;
	
`endif